`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:12:00 11/28/2018 
// Design Name: 
// Module Name:    modExp 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module modExp(
					input clk,
					input[MSGINSIZE-1:0]msgIn,
					input[KEYSIZE-1:0]key,
					input[MODSIZE-1:0]mod,
					output reg [MSGOUTSIZE-1:0]msgOut
    );
//msgOut = [msgIN^(key)] % mod

	




endmodule
